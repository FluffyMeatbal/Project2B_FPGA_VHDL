----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Remco Pieper
-- Studentnummer: 1859875
-- Create Date: 20.11.2024 19:32:54
-- Design Name: 
-- Module Name: VGA aansturing design - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package VGA_Types is                                    --array voor input registers
    type FreqArray is array(1 to 8) of std_logic_vector(1 downto 0);
end package VGA_Types;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.Numeric_STD.ALL;
use work.VGA_Types.all;

entity VGA_aansturing is
Port (
clk: in std_logic;
f: in FreqArray;
Hsync, Vsync, video_ON: out std_logic;
vgaRed, vgaGreen, vgaBlue: out std_logic_vector(3 downto 0)
);
end VGA_aansturing;

architecture Behavioral of VGA_aansturing is
signal enable: std_logic;                               --gedeelde klok 
constant prscl : integer := 4;                          --prescaler

signal xTel : integer range 0 to 1023 := 0;
signal yTel : integer range 0 to 1023 := 0;

signal H_sync : std_logic;
signal V_sync : std_logic;
signal vid_ON : std_logic;

signal Red, Green, Blue: std_logic_vector(3 downto 0);

type BlokLimiet is record
    L: integer;
    R: integer;
end record;

type BlokArray is array(1 to 8) of BlokLimiet;

constant BlokGrens: BlokArray := (                          --Array met randwaarden van de blokjes
(L => 0, R => 480/8),                                       --Blok 1
(L => 480/8+1, R => 480/8*2),                               --Blok 2
(L => 480/8*2+1, R => 480/8*3),                             --Blok 3
(L => 480/8*3+1, R => 480/8*4),                             --Blok 4
(L => 480/8*4+1, R => 480/8*5),                             --Blok 5
(L => 480/8*5+1, R => 480/8*6),                             --Blok 6
(L => 480/8*6+1, R => 480/8*7),                             --Blok 7
(L => 480/8*7+1, R => 480)                                  --Blok 8
);
constant BlockBottom:   integer := 0;                       --onderkant blokjes
constant LaagLVL:       integer := 0;                       --laag niveau blokjes
constant MediumLVL:     integer := 0;                       --medium niveau blokjes
constant HighLVL:       integer := 0;                       --hoog niveau blokjes

begin

delerBlok: process(clk)
variable deler : integer range 0 to 511 := 1;               --variabele voor de deler

begin
    if rising_edge(clk) then
        if deler = prscl / 4 then                           --25% van periode voorbij 
            enable <= '1';
        else
            enable <= '0';
        end if;
        
        if deler = prscl then                               --100% van periode voorbij 
            deler := 1;
        else
            deler := deler + 1;
        end if;
    end if;
end process delerBlok;

X_teller: process(clk, enable, xTel)
begin
    if rising_edge(clk) then
        if enable = '1' then
            if xTel < 799 then
                xTel <= xTel + 1;                           --verhoog xTel
            else
                xTel <= 0;                                  --xTel gaat terug naar het begin
            end if;
        end if;
    end if;
end process X_teller;

Y_Teller: process(clk, enable, yTel)
begin
    if rising_edge(clk) then
        if enable = '1' then
            if xTel = 799 then                              --xTel is aan het eind
                if yTel < 524 then
                    yTel <= yTel + 1;
                else 
                    yTel <= 0;
                end if;
            end if;
        end if;
    end if;
end process Y_teller;

HORsync: process(xTel)
begin
    if xTel > 655 and xTel < 752 then                       --Horizontale puls 96 lijnen breed
        H_sync <= '0';
    elsif xTel < 640 then
        H_sync <= '1';
    else
        H_sync <= '1';
    end if;
end process HORsync;

VERTsync: process(yTel)
begin
    if yTel > 489 and yTel < 492 then                       --Verticale puls 2 lijnen breed
        V_sync <= '0';
    elsif yTel < 480 then
        V_sync <= '1';
    else
        V_sync <= '1';
    end if;
end process VERTsync;

video_ON_sync: process(xTel, yTel)
begin
    if xTel < 640 and yTel < 480 then
        vid_ON <= '1';
    else
        vid_ON <= '0';
    end if;
end process video_ON_sync;

RGBsync: process(clk, enable, Red, Green, Blue, vid_ON)
begin
    if rising_edge(clk) then
        if enable = '1' then
            if vid_ON = '1' then
                vgaRed <= Red;
                vgaGreen <= Green;
                vgaBlue <= Blue;
            else
                vgaRed <= "0000";
                vgaGreen <= "0000";
                vgaBlue <= "0000";
            end if;
        end if;
    end if;
end process RGBsync;

Hsync <= H_sync;
Vsync <= V_sync;
video_ON <= vid_ON;

RegDecoder: process(clk, enable, xTel, yTel,f)

begin
    if rising_edge(clk) then
        if enable = '1' then
            for i in 1 to 8 loop                            --doorloop routine voor elke frequentie
                if xTel >= BlokGrens(i).L and xTel <= BlokGrens(i).R and yTel >= BlockBottom then  --als de x teller zich in het blokje bevind ga verder met de routine
                    if unsigned(f(i)) > 0 then
                        if yTel <= LaagLVL then             --vergelijk y teller met onderste niveau
                            Red <= "0000";                  --kleur = Groen
                            Green <= "1111";
                            Blue <= "0000";
                        end if;
                        
                        if unsigned(f(i)) > 1 then
                            if yTel <= MediumLVL then       --vergelijk y teller met middelste niveu
                                Red <= "1111";              --kleur = Geel
                                Green <= "1111";
                                Blue <= "0000";
                            end if;
                            
                            if unsigned(f(i)) > 2 then
                                if yTel <= HighLVL then     --vergelijk y teller met hoogste niveau
                                    Red <= "1111";          --kleur = Rood
                                    Green <= "0000";
                                    Blue <= "0000";
                                end if;
                            end if;
                        end if;
                    end if;
                else                                        --als de x teller niet in het blokje is dan worden de RGB signalen gelijk aan de achtergrond kleur
                    Red <= "0000";                          --achtergrond kleur = Zwart
                    Green <= "0000";
                    Blue <= "0000";
                end if;
            end loop;
        end if;
    end if;
end process RegDecoder;

end Behavioral;

